--! 
--! @file: pkg_my_data_types.vhd
--! @brief: 
--! @author: Antonio Gutierrez
--! @date: 2013-10-24
--!
--!
--------------------------------------
package my_data_types is
    type matrix is array of (natural range<>, natural range<>) of std_logic;
end package my_data_types;
------------------------------
package body my_data_types is
    --functionsdefinitions
end package body my_data_types;
--------------------------------------

