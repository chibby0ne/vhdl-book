------------------------------
package my_data_type is 
    type oneDoneD is array (0 to 3) of bit_vector(7 downto 0);
end package;
------------------------------

