--! 
--! @file: exercise6_13.vhd
--! @brief: Programmable signal generator with frequency meter
--! @author: Antonio Gutierrez
--! @date: 2013-10-28
--!
--!
--------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_all;
--------------------------------------
entity program_signal_generator_with_freq_meter is
--generic declarations
    port (
        in: in std_logic;
        out: out std_logic);
end entity program_signal_generator_with_freq_meter;
--------------------------------------
architecture circuit of program_signal_generator_with_freq_meter is
--signals and declarations
begin
    --architecture_statements_part
end architecture circuit;

